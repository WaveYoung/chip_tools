`ifndef BENCH_PKG_SV
`define BENCH_PKG_SV

//common_lib
`include "common_lib/lib_pkg.sv"

//include package file

//import packages

//include files
`include "virtual_sequencer.sv"
`include "virtual_sequence.sv"
`include "base_test.sv"
`include "assert/examp_assert.sv"
`include "tb_top.sv"

`endif