`ifndef TESTCASE_PKG_SV
`define TESTCASE_PKG_SV

//include package file

//import packages

//include files
`include "example_case.sv"

`endif