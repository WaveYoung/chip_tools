`ifndef LIB_PKG_SV
`define LIB_PKG_SV

// import uvm package
import uvm_pkg::*;
`include "uvm_macros.svh"
// include common lib module
`include "clk_gen.sv"
`include "dump_wave.sv"

`endif
